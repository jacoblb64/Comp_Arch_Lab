--library ieee;
--use ieee.std_logic_1164.all; -- allows use of the std_logic_vector type
----use ieee.std_logic_arith.all;
----use ieee.std_logic_unsigned.all;
--use ieee.numeric_std.all;

--entity ALU_tb is
--end entity ; -- ALU_tb

--architecture arch of ALU_tb is
	
--	component ALU_tb is
--	  port (
--		clock
--	  ) ;
--	end component ; -- ALU_tb


--begin



--end architecture ; -- arch