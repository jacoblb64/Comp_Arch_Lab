--library ieee;
--use ieee.std_logic_1164.all; -- allows use of the std_logic_vector type
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--use ieee.numeric_std.all;
--
--library lpm;
--use lpm.lpm_components.all;
--
--entity key_inverter is
--
--end key_inverter;
--
--architecture struct of key_inverter is
--
--	signal 
--
--begin
--
--end architecture ; -- struct