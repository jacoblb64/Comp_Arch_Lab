library verilog;
use verilog.vl_types.all;
entity matrix_multiplier_vlg_vec_tst is
end matrix_multiplier_vlg_vec_tst;
